module gold_mult(
input clk,
input reset_n,
input [15:0] a,
input [15:0] b,
output [31:0] result
);
// TODO: Implement the multiplication of a and b and store the result in result
// This should be the reference implementation that we compare test_mult against

endmodule