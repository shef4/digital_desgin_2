`ifndef STATUS_DEFS_SV
`define STATUS_DEFS_SV

`timescale 1ns/1ns
`default_nettype none




`endif // STATUS_DEFS_SV