// audio_fifo.v

// Generated using ACDS version 22.1 915

`timescale 1 ps / 1 ps
module audio_fifo (
		input  wire        sc_fifo_0_clk_clk,         //       sc_fifo_0_clk.clk
		input  wire        sc_fifo_0_clk_reset_reset, // sc_fifo_0_clk_reset.reset
		input  wire [15:0] sc_fifo_0_in_data,         //        sc_fifo_0_in.data
		input  wire        sc_fifo_0_in_valid,        //                    .valid
		output wire        sc_fifo_0_in_ready,        //                    .ready
		output wire [15:0] sc_fifo_0_out_data,        //       sc_fifo_0_out.data
		output wire        sc_fifo_0_out_valid,       //                    .valid
		input  wire        sc_fifo_0_out_ready        //                    .ready
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (16),
		.FIFO_DEPTH          (1024),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (0),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (3),
		.USE_MEMORY_BLOCKS   (1),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) sc_fifo_0 (
		.clk               (sc_fifo_0_clk_clk),                    //       clk.clk
		.reset             (sc_fifo_0_clk_reset_reset),            // clk_reset.reset
		.in_data           (sc_fifo_0_in_data),                    //        in.data
		.in_valid          (sc_fifo_0_in_valid),                   //          .valid
		.in_ready          (sc_fifo_0_in_ready),                   //          .ready
		.out_data          (sc_fifo_0_out_data),                   //       out.data
		.out_valid         (sc_fifo_0_out_valid),                  //          .valid
		.out_ready         (sc_fifo_0_out_ready),                  //          .ready
		.csr_address       (2'b00),                                // (terminated)
		.csr_read          (1'b0),                                 // (terminated)
		.csr_write         (1'b0),                                 // (terminated)
		.csr_readdata      (),                                     // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000), // (terminated)
		.almost_full_data  (),                                     // (terminated)
		.almost_empty_data (),                                     // (terminated)
		.in_startofpacket  (1'b0),                                 // (terminated)
		.in_endofpacket    (1'b0),                                 // (terminated)
		.out_startofpacket (),                                     // (terminated)
		.out_endofpacket   (),                                     // (terminated)
		.in_empty          (1'b0),                                 // (terminated)
		.out_empty         (),                                     // (terminated)
		.in_error          (1'b0),                                 // (terminated)
		.out_error         (),                                     // (terminated)
		.in_channel        (1'b0),                                 // (terminated)
		.out_channel       ()                                      // (terminated)
	);

endmodule
