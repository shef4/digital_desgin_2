

module mult16_tester(
    input         CLOCK_50, 
    input  [2:0]  KEY, 
    output [6:0]  HEX5, 
    output [6:0]  HEX4,
    output [6:0]  HEX3, 
    output [6:0]  HEX2, 
    output [6:0]  HEX1, 
    output [6:0]  HEX0
);

    reg 			 clock;
    wire [31:0] test_result, gold_result;
    wire        match,busy, begin_test, inject_error;
    wire        test_mult_start;
	logic 		reset;
	logic [1:0] reset_int;
	logic [4:0] status_out;
	logic [15:0] opA, opB;
    

    
    // button debouncing and edge detection
	// Define the first flip-flop stage
	always_ff @(posedge CLOCK_50)
		reset_int[0] <= KEY[0];

	// Define the second flip-flop stage
	always_ff @(posedge CLOCK_50)
		reset_int[1] <= reset_int[0];

	// Define the output flip-flop stage
	always_ff @(posedge CLOCK_50)
		reset <= reset_int[1];
		
	// clock divider to generate 1Hz clock
	always @(posedge CLOCK_50) begin
        if (!reset) begin
            clock <= 0;
        end else if (clock) begin
            clock <= 0;
        end else begin
            clock <= 1;
        end
   end

											
	button start_debounce(  .clock(clock), 
							.reset(reset), 
							.button_in(KEY[1]), 
							.pulse_out(begin_test));
											
	button error_debounce( 	.clock(clock), 
							.reset(reset), 
							.button_in(KEY[1]), 
							.pulse_out(inject_error));
    
    // status module to output the status register to the HEX displays
    status status_inst(	.clock(CLOCK_50), .reset_n(reset),
					   	.begin_test(begin_test), .inject_error(inject_error),
					   	.busy(busy),.results_match(match),
						.status_out(status_out), 
						.opA(opA), .opB(opB),
						.test_mult_start(test_mult_start));
							  
    // test multiplier to calculate product of A and B
    test_mult test_mult_inst(.clk(clock),.reset_n(reset),.start(test_mult_start),
							.a(opA), .b(opB),
							.busy(busy),.result(test_result));
    
    // gold standard multiplier to calculate product of A and B
    gold_mult gold_mult_inst(.a(opA),.b(opB),.result(gold_result));
    
    // comparator to check if the test multiplier matches the gold multiplier
    compare compare_inst(.test_result(test_result), .gold_result(gold_result),.match(match));
    
    // output the status register to the HEX displays
	seg_disp seg_disp_inst5(.clock(clock),.num(status_out),.seg(HEX5));
	seg_disp seg_disp_inst4(.clock(clock),.num(status_out),.seg(HEX4));
	seg_disp seg_disp_inst3(.clock(clock),.num({1'b0,opA[15:12]}),.seg(HEX3));
	seg_disp seg_disp_inst2(.clock(clock),.num({1'b0,opA[11:8]}),.seg(HEX2));
	seg_disp seg_disp_inst1(.clock(clock),.num({1'b0,opB[15:12]}),.seg(HEX1));
	seg_disp seg_disp_inst0(.clock(clock),.num({1'b0,opB[11:8]}),.seg(HEX0));
		  
endmodule

module mult16_tester_tb;
	// Inputs
	reg         CLOCK_50;
	reg  [2:0]  KEY;

	// Outputs
	wire [6:0]  HEX5;
	wire [6:0]  HEX4;
	wire [6:0]  HEX3;
	wire [6:0]  HEX2;
	wire [6:0]  HEX1;
	wire [6:0]  HEX0;

	// Instantiate the Unit Under Test (UUT)
	mult16_tester uut (
		 .CLOCK_50(CLOCK_50), 
		 .KEY(KEY), 
		 .HEX5(HEX5), 
		 .HEX4(HEX4), 
		 .HEX3(HEX3), 
		 .HEX2(HEX2), 
		 .HEX1(HEX1), 
		 .HEX0(HEX0)
	);

	initial begin
		 // Initialize Inputs
		 CLOCK_50 = 0;
		 KEY = 0;

		 // Wait 100 ns for global reset to finish
		 #100;

		 // Add stimulus here
		 KEY = 1; // Press the start button
		 #100;
		 KEY = 0; // Release the start button
		 #20000;

		 $finish;
	end

	always #25 CLOCK_50 = ~CLOCK_50;
endmodule
