`ifndef MULT16_TESTER_DEFS_SV
`define MULT16_TESTER_DEFS_SV

`timescale 1ns/1ps
`default_nettype none


// Define user-defined data types
// TODO: Add any user-defined data types required in multiple source files

`endif // MULT16_TESTER_DEFS_SV