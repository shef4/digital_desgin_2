module test_mult(
input clk,
input reset_n,
input [15:0] a,
input [15:0] b,
output [31:0] result
);
// TODO: Add your code here
endmodule