`ifndef MULT16_TESTER_DEFS_SV
`define MULT16_TESTER_DEFS_SV





`endif
