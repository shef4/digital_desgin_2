// audio_controller.v

// Generated using ACDS version 22.1 915

`timescale 1 ps / 1 ps
module audio_controller (
		input  wire [15:0] audio_0_avalon_left_channel_sink_data,   //  audio_0_avalon_left_channel_sink.data
		input  wire        audio_0_avalon_left_channel_sink_valid,  //                                  .valid
		output wire        audio_0_avalon_left_channel_sink_ready,  //                                  .ready
		input  wire [15:0] audio_0_avalon_right_channel_sink_data,  // audio_0_avalon_right_channel_sink.data
		input  wire        audio_0_avalon_right_channel_sink_valid, //                                  .valid
		output wire        audio_0_avalon_right_channel_sink_ready, //                                  .ready
		input  wire        audio_0_clk_clk,                         //                       audio_0_clk.clk
		input  wire        audio_0_external_interface_BCLK,         //        audio_0_external_interface.BCLK
		output wire        audio_0_external_interface_DACDAT,       //                                  .DACDAT
		input  wire        audio_0_external_interface_DACLRCK,      //                                  .DACLRCK
		input  wire        audio_0_reset_reset                      //                     audio_0_reset.reset
	);

	audio_controller_audio_0 audio_0 (
		.clk                          (audio_0_clk_clk),                         //                         clk.clk
		.reset                        (audio_0_reset_reset),                     //                       reset.reset
		.from_adc_left_channel_ready  (),                                        //  avalon_left_channel_source.ready
		.from_adc_left_channel_data   (),                                        //                            .data
		.from_adc_left_channel_valid  (),                                        //                            .valid
		.from_adc_right_channel_ready (),                                        // avalon_right_channel_source.ready
		.from_adc_right_channel_data  (),                                        //                            .data
		.from_adc_right_channel_valid (),                                        //                            .valid
		.to_dac_left_channel_data     (audio_0_avalon_left_channel_sink_data),   //    avalon_left_channel_sink.data
		.to_dac_left_channel_valid    (audio_0_avalon_left_channel_sink_valid),  //                            .valid
		.to_dac_left_channel_ready    (audio_0_avalon_left_channel_sink_ready),  //                            .ready
		.to_dac_right_channel_data    (audio_0_avalon_right_channel_sink_data),  //   avalon_right_channel_sink.data
		.to_dac_right_channel_valid   (audio_0_avalon_right_channel_sink_valid), //                            .valid
		.to_dac_right_channel_ready   (audio_0_avalon_right_channel_sink_ready), //                            .ready
		.AUD_BCLK                     (audio_0_external_interface_BCLK),         //          external_interface.export
		.AUD_DACDAT                   (audio_0_external_interface_DACDAT),       //                            .export
		.AUD_DACLRCK                  (audio_0_external_interface_DACLRCK)       //                            .export
	);

endmodule
