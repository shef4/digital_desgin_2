module compare(
input clk,
input reset_n,
input [31:0] test_mult,
input [31:0] gold_mult,
output match
);

endmodule